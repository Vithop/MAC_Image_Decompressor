library verilog;
use verilog.vl_types.all;
entity Milestone1_v_unit is
end Milestone1_v_unit;
