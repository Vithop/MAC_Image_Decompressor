library verilog;
use verilog.vl_types.all;
entity MAC_Image_Decompressor_v_unit is
end MAC_Image_Decompressor_v_unit;
