
`timescale 1ns/100ps

`ifndef DISABLE_DEFAULT_NET
`default_nettype none
`endif

module multiplier (	
	output logic [31:0] a
	input logic [31:0] b,
	input logic [31:0] c,
	
	output logic [31:0] d,
	input logic [31:0] e,
	input logic [31:0] f,

	output logic [31:0] g,
	input logic [31:0] h,
	input logic [31:0] i,
);

	
endmodule
