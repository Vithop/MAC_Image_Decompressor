
`timescale 1ns/100ps

`ifndef DISABLE_DEFAULT_NET
`default_nettype none
`endif

module multiplier (
	input logic [31:0] a,
	input logic [31:0] b,
	output logic [63:0] c
);

always_comb begin
	case()
		
	endcase
end
	
endmodule
